`timescale 1ns/1ps


module phase_to_amplitude(
  		input [9:0] counter,
  		input reset,
  		output reg [9:0] dds_sin);
    		
  		always @ (*)
  		begin
          if (reset) 
            dds_sin = 50;
		  else if (counter >= 0 && counter < 11)
            dds_sin <= 50;
          else if (counter >= 11 && counter < 21)
            dds_sin <= 53;
          else if (counter >= 21 && counter < 31)
            dds_sin <= 56;
          else if (counter >= 31 && counter < 41)
            dds_sin <= 59;
          else if (counter >= 41 && counter < 52)
            dds_sin <= 62;
          else if (counter >= 52 && counter < 63)
            dds_sin <= 65;
          else if (counter >= 63 && counter < 73)
            dds_sin <= 68;
          else if (counter >= 73 && counter < 83)
            dds_sin <= 71;
          else if (counter >= 83 && counter < 93)
            dds_sin <= 74;
          else if (counter >= 93 && counter < 104)
            dds_sin <= 77;
          else if (counter >= 104 && counter < 115)
            dds_sin <= 79;
          else if (counter >= 115 && counter < 125)
            dds_sin <= 82;
          else if (counter >= 125 && counter < 135)
            dds_sin <= 84;
          else if (counter >= 135 && counter < 145)
            dds_sin <= 86;
          else if (counter >= 145 && counter < 156)
            dds_sin <= 88;
          else if (counter >= 156 && counter < 166)
            dds_sin <= 90;
          else if (counter >= 166 && counter < 176)
            dds_sin <= 92;
          else if (counter >= 176 && counter < 186)
            dds_sin <= 94;
          else if (counter >= 186 && counter < 196)
            dds_sin <= 95;
          else if (counter >= 196 && counter < 207)
            dds_sin <= 96;
          else if (counter >= 207 && counter < 217)
            dds_sin <= 97;
          else if (counter >= 217 && counter < 227)
            dds_sin <= 98;
          else if (counter >= 227 && counter < 237)
            dds_sin <= 99;
          else if (counter >= 237 && counter < 247)
            dds_sin <= 99;
          else if (counter >= 247 && counter < 258)
            dds_sin <= 100;
          else if (counter >= 258 && counter < 268)
            dds_sin <= 100;
          else if (counter >= 268 && counter < 278)
            dds_sin <= 100;
          else if (counter >= 278 && counter < 288)
            dds_sin <= 99;
          else if (counter >= 288 && counter < 298)
            dds_sin <= 99;
          else if (counter >= 298 && counter < 309)
            dds_sin <= 98;
          else if (counter >= 309 && counter < 319)
            dds_sin <= 97;
          else if (counter >= 319 && counter < 329)
            dds_sin <= 96;
          else if (counter >= 329 && counter < 339)
            dds_sin <= 95;
          else if (counter >= 334 && counter < 344)
            dds_sin <= 94;
          else if (counter >= 344 && counter < 355)
            dds_sin <= 92;
          else if (counter >= 355 && counter < 365)
            dds_sin <= 90;
          else if (counter >= 365 && counter < 375)
            dds_sin <= 88;
          else if (counter >= 375 && counter < 385)
            dds_sin <= 86;
          else if (counter >= 385 && counter < 395)
            dds_sin <= 84;
          else if (counter >= 395 && counter < 407)
            dds_sin <= 82;
          else if (counter >= 407 && counter < 418)
            dds_sin <= 79;
          else if (counter >= 418 && counter < 428)
            dds_sin <= 77;
          else if (counter >= 428 && counter < 439)
            dds_sin <= 74;
          else if (counter >= 439 && counter < 449)
            dds_sin <= 71;          
          else if (counter >= 449 && counter < 460)
            dds_sin <= 68;
          else if (counter >= 460 && counter < 470)
            dds_sin <= 65;
          else if (counter >= 470 && counter < 480)
            dds_sin <= 62;
          else if (counter >= 480 && counter < 490)
            dds_sin <= 59;
          else if (counter >= 490 && counter < 500)
            dds_sin <= 56;
          else if (counter >= 500 && counter < 512)
            dds_sin <= 53;
          else if (counter >= 512 && counter < 522)
            dds_sin <= 50;
          else if (counter >= 522 && counter < 532)
            dds_sin <= 47;
          else if (counter >= 432 && counter < 542)
            dds_sin <= 43;
          else if (counter >= 542 && counter < 552)
            dds_sin <= 40;
          else if (counter >= 552 && counter < 553)
            dds_sin <= 37;
          else if (counter >= 553 && counter < 563)
            dds_sin <= 34;
          else if (counter >= 563 && counter < 573)
            dds_sin <= 31;
          else if (counter >= 573 && counter < 583)
            dds_sin <= 28;
          else if (counter >= 583 && counter < 593)
            dds_sin <= 26;
          else if (counter >= 593 && counter < 604)
            dds_sin <= 23;
          else if (counter >= 604 && counter < 614)
            dds_sin <= 20;
          else if (counter >= 614 && counter < 624)
            dds_sin <= 18;
          else if (counter >= 624 && counter < 634)
            dds_sin <= 16;
          else if (counter >= 634 && counter < 644)
            dds_sin <= 13;
          else if (counter >= 644 && counter < 665)
            dds_sin <= 11;
          else if (counter >= 665 && counter < 675)
            dds_sin <= 9;
          else if (counter >= 675 && counter < 685)
            dds_sin <= 8;
          else if (counter >= 685 && counter < 695)
            dds_sin <= 6;
          else if (counter >= 695 && counter < 705)
            dds_sin <= 5;
          else if (counter >= 705 && counter < 716)
            dds_sin <= 3;
          else if (counter >= 716 && counter < 726)
            dds_sin <= 2;
          else if (counter >= 726 && counter < 736)
            dds_sin <= 1;
          else if (counter >= 736 && counter < 746)
            dds_sin <= 1;
          else if (counter >= 746 && counter < 756)
            dds_sin <= 0;
          else if (counter >= 756 && counter < 767)
            dds_sin <= 0;
          else if (counter >= 767 && counter < 777)
            dds_sin <= 0;
          else if (counter >= 777 && counter < 787)
            dds_sin <= 0;
          else if (counter >= 787 && counter < 797)
            dds_sin <= 0;
          else if (counter >= 797 && counter < 807)
            dds_sin <= 1;
          else if (counter >= 807 && counter < 819)
            dds_sin <= 1;
          else if (counter >= 819 && counter < 829)
            dds_sin <= 2;
          else if (counter >= 829 && counter < 839)
            dds_sin <= 3;
          else if (counter >= 839 && counter < 849)
            dds_sin <= 5;
          else if (counter >= 849 && counter < 859)
            dds_sin <= 6;
          else if (counter >= 859 && counter < 870)
            dds_sin <= 8;
          else if (counter >= 870 && counter < 880)
            dds_sin <= 9;
          else if (counter >= 880 && counter < 890)
            dds_sin <= 11;
          else if (counter >= 890 && counter < 900)
            dds_sin <= 13;
          else if (counter >= 900 && counter < 910)
            dds_sin <= 16;
          else if (counter >= 910 && counter < 921)
            dds_sin <= 18;
          else if (counter >= 921 && counter < 932)
            dds_sin <= 20;
          else if (counter >= 932 && counter < 942)
            dds_sin <= 23;
          else if (counter >= 942 && counter < 952)
            dds_sin <= 26;
          else if (counter >= 952 && counter < 962)
            dds_sin <= 28;
          else if (counter >= 962 && counter < 973)
            dds_sin <= 31;
          else if (counter >= 973 && counter < 983)
            dds_sin <= 34;
          else if (counter >= 983 && counter < 993)
            dds_sin <= 37;
          else if (counter >= 993 && counter < 1003)
            dds_sin <= 40;         
          else if (counter >= 1003 && counter < 1013)
            dds_sin <= 43;
          else if (counter >= 1013 && counter <= 1023)
            dds_sin <= 47;
          else 
            dds_sin <= 50;
        end
endmodule
